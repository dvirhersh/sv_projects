`ifndef CFS_ALGN_ENV_SV
	`define CFS_ALGN_ENV_SV

	class cfs_algn_env extends uvm_env;
		
	endclass : cfs_algn_env

`endif