`ifndef CFS_APB_PKG_SV
	`define CFS_APB_PKG_SV

	`include "uvm_macros.svh"

	package cfs_apb_pkg;
		import uvm_pkg::*;

	endpackage

`endif