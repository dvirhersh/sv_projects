class pmulticast extends packet;
  function new(input string name = "pmulticast");
    super.new();
  endfunction
endclass
