class psingle extends packet;
  function new(input string name = "psingle");
    super.new();
  endfunction
endclass
