class psingle extends packet;
    function new(input string name = "psingle");
        super.new(name);
    endfunction
endclass
